library ieee;
use ieee.std_logic_1164.all;

entity mux2to1 is
port
	(
		d0		:	in 	std_logic_vector(3 downto 0);
		d1		:	in		std_logic_vector(3 downto 0);
		d2		:	in		std_logic_vector(3 downto 0);
		d3		:	in		std_logic_vector(3 downto 0);
		s		:	in		std_logic_vector(1 downto 0);
		F		:	out	std_logic_vector(3 downto 0)
	);
end mux2to1;

architecture logicFunction of mux2to1 is

begin
	with s select
		f <= 	d0 when "00",
				d1 when "01",
				d2 when "10",
				d3 when "11";
end logicFunction;